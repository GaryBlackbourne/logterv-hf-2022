`timescale 1ns / 1ps

module top(
    input clk,
    input rst
    
    // todo: FPGA lábak és CODEC jelek
    
    );
    
    codec_if codec_interface(
        // todo: wiring
    );
    
    flanger flanger_effect(
        // todo: wiring
    );
    
endmodule
